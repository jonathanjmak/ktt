//
//  music_player module
//
//  This music_player module connects up the MCU, song_reader, note_player,
//  beat_generator, and codec_conditioner. It provides an output that indicates
//  a new sample (new_sample_generated) which will be used in lab 5.
//

module music_player(
    // Standard system clock and reset
    input clk,
    input reset,

    // Our debounced and one-pulsed button inputs.
    input play_button,
    input next_button,

    // The raw  signal from the ac97_if codec.
    input new_frame,

    // This output must go high for one cycle when a new sample is generated.
    output wire new_sample_generated,

    // Our final output sample to the codec. This needs to be synced to
    // new_frame.
    output wire [15:0] sample_out
);
    // The BEAT_COUNT is parameterized so you can reduce this in simulation.
    // If you reduce this to 100 your simulation will be 10x faster.
    parameter BEAT_COUNT = 1000;


//
//  ****************************************************************************
//      Master Control Unit
//  ****************************************************************************
//   The reset_player output from the MCU is run only to the song_reader because
//   we don't need to reset any state in the note_player. If we do it may make
//   a pop when it resets the output sample.
//
 
    wire play;
    wire reset_player;
    wire [1:0] current_song;
    wire song_done;
    mcu mcu(
        .clk(clk),
        .reset(reset),
        .play_button(play_button),
        .next_button(next_button),
        .play(play),
        .reset_player(reset_player),
        .song(current_song),
        .song_done(song_done)
    );
	 

//
//  ****************************************************************************
//      Song Reader
//  ****************************************************************************
//
    wire [5:0] note_to_play;
    wire [5:0] duration_for_note;
    wire new_note;
	 wire player_ready;
	 wire beat;

//	song_reader song_reader(
//		.clk(clk),
//		.reset(reset | reset_player),
//		.play(play),
//		.player_ready(player_ready),
//		.song(current_song),
//		.beat(beat),
//		.song_done(song_done),
//		.note(note_to_play),
//		.duration(duration_for_note),
//		.new_note(new_note)
//   );

		song_reader song_reader(
		.clk(clk),
		.reset(reset | reset_player),
		.play(play),
		.player_available(player_ready),
		.song(current_song),
		.beat(beat),
		.song_done(song_done),
		.note(note_to_play),
		.duration(duration_for_note),
		.new_note(new_note)
   );
//
//  ****************************************************************************
//      Chords Module
//  ****************************************************************************
//
		wire generate_next_sample;
		wire [15:0] note_sample;
		wire note_sample_ready;
	 
		chords chord_module(	
			.clk(clk), 
			.reset(reset|reset_player),
			.play(play),
			.note(note_to_play),
			.duration(duration_for_note),
			.new_note(new_note),
			.beat(beat),
			.generate_next_sample(generate_next_sample),
			.player_ready(player_ready),
			.sample_out(note_sample),
			.new_sample_ready(note_sample_ready)
		);
      
//   
//  ****************************************************************************
//      Beat Generator
//  ****************************************************************************
//  By default this will divide the generate_next_sample signal (48kHz from the
//  codec's new_frame input) down by 1000, to 48Hz. If you change the BEAT_COUNT
//  parameter when instantiating this you can change it for simulation.
//  
    beat_generator #(.WIDTH(10), .STOP(BEAT_COUNT)) beat_generator(
        .clk(clk),
        .reset(reset),
        .en(generate_next_sample),
        .beat(beat)
    );

//  
//  ****************************************************************************
//      Codec Conditioner
//  ****************************************************************************
//  
    assign new_sample_generated = generate_next_sample;
    codec_conditioner codec_conditioner(
        .clk(clk),
        .reset(reset),
        .new_sample_in(note_sample),
        .latch_new_sample_in(note_sample_ready),
        .generate_next_sample(generate_next_sample),
        .new_frame(new_frame),
        .valid_sample(sample_out)
    );

endmodule
