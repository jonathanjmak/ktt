// // How to use:					
// // 1. Edit the songs on the Enter Song sheet.					
// // 2. Select this whole worksheet, copy it, and paste it into a new file.					
// // 3. Save the file as song_rom.v.					
					
// // A test song_rom with the new song format. 				
// module song_rom (					
// 	input clk,				
// 	input [10:0] addr,				
// 	output reg [15:0] dout				
// );					
					
// 	wire [15:0] memory [2047:0];				
					
// 	always @(posedge clk)				
// 		dout = memory[addr];			
					
// 	assign memory[	  0	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	  1	] =	{1'b0,6'd32, 6'd12,3'b111};	// Note: 3E
// 	assign memory[	  2	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	  3	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	  4	] =	{1'b0,6'd33, 6'd12,3'b111};	// Note: 3F
// 	assign memory[	  5	] =	{1'b0,6'd37, 6'd12,3'b111};	// Note: 4A
// 	assign memory[	  6	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	  7	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	  8	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	  9	] =	{1'b0,6'd39, 6'd12,3'b111};	// Note: 4B
// 	assign memory[	 10	] =	{1'b0,6'd42, 6'd12,3'b111};	// Note: 4D
// 	assign memory[	 11	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 12	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 13	] =	{1'b0,6'd44, 6'd12,3'b111};	// Note: 4E
// 	assign memory[	 14	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 15	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 16	] =	{1'b0,6'd45, 6'd12,3'b111};	// Note: 4F
// 	assign memory[	 17	] =	{1'b0,6'd49, 6'd12,3'b111};	// Note: 5A
// 	assign memory[	 18	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 19	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 20	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 21	] =	{1'b0,6'd51, 6'd12,3'b111};	// Note: 5B
// 	assign memory[	 22	] =	{1'b0,6'd54, 6'd12,3'b111};	// Note: 5D
// 	assign memory[	 23	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 24	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 25	] =	{1'b0,6'd55, 6'd12,3'b111};	// Note: 5D#Eb
// 	assign memory[	 26	] =	{1'b0,6'd58, 6'd12,3'b111};	// Note: 5F#Gb
// 	assign memory[	 27	] =	{1'b0,6'd0, 6'd12,3'b111};	// Note: rest
// 	assign memory[	 28	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 29	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 30	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 31	] =	{1'b1,6'd0, 6'd0,3'b111};	// Note: rest
// 	assign memory[	 32	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 33	] =	{1'b0,6'd32, 6'd12,3'b111};	// Note: 3E
// 	assign memory[	 34	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	 35	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 36	] =	{1'b0,6'd33, 6'd12,3'b111};	// Note: 3F
// 	assign memory[	 37	] =	{1'b0,6'd37, 6'd12,3'b111};	// Note: 4A
// 	assign memory[	 38	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 39	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 40	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	 41	] =	{1'b0,6'd39, 6'd12,3'b111};	// Note: 4B
// 	assign memory[	 42	] =	{1'b0,6'd42, 6'd12,3'b111};	// Note: 4D
// 	assign memory[	 43	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 44	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 45	] =	{1'b0,6'd44, 6'd12,3'b111};	// Note: 4E
// 	assign memory[	 46	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 47	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 48	] =	{1'b0,6'd45, 6'd12,3'b111};	// Note: 4F
// 	assign memory[	 49	] =	{1'b0,6'd49, 6'd12,3'b111};	// Note: 5A
// 	assign memory[	 50	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 51	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 52	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 53	] =	{1'b0,6'd51, 6'd12,3'b111};	// Note: 5B
// 	assign memory[	 54	] =	{1'b0,6'd54, 6'd12,3'b111};	// Note: 5D
// 	assign memory[	 55	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 56	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 57	] =	{1'b0,6'd55, 6'd12,3'b111};	// Note: 5D#Eb
// 	assign memory[	 58	] =	{1'b0,6'd58, 6'd12,3'b111};	// Note: 5F#Gb
// 	assign memory[	 59	] =	{1'b0,6'd0, 6'd12,3'b111};	// Note: rest
// 	assign memory[	 60	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 61	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 62	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 63	] =	{1'b1,6'd0, 6'd0,3'b111};	// Note: rest
// 	assign memory[	 64	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 65	] =	{1'b0,6'd32, 6'd12,3'b111};	// Note: 3E
// 	assign memory[	 66	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	 67	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 68	] =	{1'b0,6'd33, 6'd12,3'b111};	// Note: 3F
// 	assign memory[	 69	] =	{1'b0,6'd37, 6'd12,3'b111};	// Note: 4A
// 	assign memory[	 70	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 71	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 72	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	 73	] =	{1'b0,6'd39, 6'd12,3'b111};	// Note: 4B
// 	assign memory[	 74	] =	{1'b0,6'd42, 6'd12,3'b111};	// Note: 4D
// 	assign memory[	 75	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 76	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 77	] =	{1'b0,6'd44, 6'd12,3'b111};	// Note: 4E
// 	assign memory[	 78	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 79	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 80	] =	{1'b0,6'd45, 6'd12,3'b111};	// Note: 4F
// 	assign memory[	 81	] =	{1'b0,6'd49, 6'd12,3'b111};	// Note: 5A
// 	assign memory[	 82	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 83	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 84	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	 85	] =	{1'b0,6'd51, 6'd12,3'b111};	// Note: 5B
// 	assign memory[	 86	] =	{1'b0,6'd54, 6'd12,3'b111};	// Note: 5D
// 	assign memory[	 87	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	 88	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 89	] =	{1'b0,6'd55, 6'd12,3'b111};	// Note: 5D#Eb
// 	assign memory[	 90	] =	{1'b0,6'd58, 6'd12,3'b111};	// Note: 5F#Gb
// 	assign memory[	 91	] =	{1'b0,6'd0, 6'd12,3'b111};	// Note: rest
// 	assign memory[	 92	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 93	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	 94	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	 95	] =	{1'b1,6'd0, 6'd0,3'b111};	// Note: rest
// 	assign memory[	 96	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	 97	] =	{1'b0,6'd32, 6'd12,3'b111};	// Note: 3E
// 	assign memory[	 98	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	 99	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	100	] =	{1'b0,6'd33, 6'd12,3'b111};	// Note: 3F
// 	assign memory[	101	] =	{1'b0,6'd37, 6'd12,3'b111};	// Note: 4A
// 	assign memory[	102	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	103	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	104	] =	{1'b0,6'd35, 6'd12,3'b111};	// Note: 3G
// 	assign memory[	105	] =	{1'b0,6'd39, 6'd12,3'b111};	// Note: 4B
// 	assign memory[	106	] =	{1'b0,6'd42, 6'd12,3'b111};	// Note: 4D
// 	assign memory[	107	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	108	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	109	] =	{1'b0,6'd44, 6'd12,3'b111};	// Note: 4E
// 	assign memory[	110	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	111	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	112	] =	{1'b0,6'd45, 6'd12,3'b111};	// Note: 4F
// 	assign memory[	113	] =	{1'b0,6'd49, 6'd12,3'b111};	// Note: 5A
// 	assign memory[	114	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	115	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	116	] =	{1'b0,6'd47, 6'd12,3'b111};	// Note: 4G
// 	assign memory[	117	] =	{1'b0,6'd51, 6'd12,3'b111};	// Note: 5B
// 	assign memory[	118	] =	{1'b0,6'd54, 6'd12,3'b111};	// Note: 5D
// 	assign memory[	119	] =	{1'b1,6'd0, 6'd8,3'b111};	// Note: rest
// 	assign memory[	120	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	121	] =	{1'b0,6'd55, 6'd12,3'b111};	// Note: 5D#Eb
// 	assign memory[	122	] =	{1'b0,6'd58, 6'd12,3'b111};	// Note: 5F#Gb
// 	assign memory[	123	] =	{1'b0,6'd0, 6'd12,3'b111};	// Note: rest
// 	assign memory[	124	] =	{1'b0,6'd28, 6'd12,3'b111};	// Note: 3C
// 	assign memory[	125	] =	{1'b0,6'd40, 6'd12,3'b111};	// Note: 4C
// 	assign memory[	126	] =	{1'b0,6'd52, 6'd12,3'b111};	// Note: 5C
// 	assign memory[	127	] =	{1'b1,6'd0, 6'd0,3'b111};	// Note: rest

// endmodule					

// A test song_rom with the new song format. 				
module song_rom (					
	input clk,				
	input [10:0] addr,				
	output reg [15:0] dout				
);					
					
	wire [15:0] memory [2047:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
	assign memory[	  0	] =	{1'b0, 6'd30, 6'd48, 3'b111};	// Note: 3D
	assign memory[	  1	] =	{1'b0, 6'd38, 6'd48, 3'b111};	// Note: 4A#Bb
	assign memory[	  2	] =	{1'b0, 6'd14, 6'd24, 3'b111};	// Note: 2A#Bb
	assign memory[	  3	] =	{1'b1, 6'd00, 6'd24, 3'b111};	// Note: rest

	assign memory[	  4	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	  5	] =	{1'b1, 6'd00, 6'd8, 3'b111};	// Note: rest
	
	assign memory[	  6	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	  7	] =	{1'b1, 6'd0, 6'd00, 3'b111};	// Note: rest (for 0)
	assign memory[	  8	] =	{1'b1, 6'd0, 6'd08, 3'b111};	// Note: rest
	
	assign memory[	  9	] =	{1'b0, 6'd14, 6'd24, 3'b111};	// Note: 2A#Bb
	assign memory[	 10	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	 11	] =	{1'b0, 6'd30, 6'd6, 3'b111};	// Note: 3D
	assign memory[	 12	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	 13	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 14	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	 15	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 16	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	 17	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 18	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	 19	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 20	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	 21	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 22	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	 23	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 24	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	 25	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 26	] =	{1'b0, 6'd38, 6'd18, 3'b111};	// Note: 4A#Bb
	assign memory[	 27	] =	{1'b0, 6'd28, 6'd18, 3'b111};	// Note: 3C
	assign memory[	 28	] =	{1'b0, 6'd12, 6'd24, 3'b111};	// Note: 1G#Ab
	assign memory[	 29	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	 30	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	 31	] =	{1'b0, 6'd28, 6'd6, 3'b111};	// Note: 3C
	assign memory[	 32	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 33	] =	{1'b0, 6'd38, 6'd36, 3'b111};	// Note: 4A#Bb
	assign memory[	 34	] =	{1'b0, 6'd28, 6'd48, 3'b111};	// Note: 3C
	assign memory[	 35	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 36	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 37	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 38	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 39	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 40	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 41	] =	{1'b0, 6'd12, 6'd24, 3'b111};	// Note: 1G#Ab
	assign memory[	 42	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	 43	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	 44	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 45	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	 46	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 47	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 48	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 49	] =	{1'b0, 6'd28, 6'd8, 3'b111};	// Note: 3C
	assign memory[	 50	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 51	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 52	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 53	] =	{1'b0, 6'd28, 6'd8, 3'b111};	// Note: 3C
	assign memory[	 54	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 55	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 56	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	 57	] =	{1'b0, 6'd28, 6'd8, 3'b111};	// Note: 3C
	assign memory[	 58	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 59	] =	{1'b0, 6'd38, 6'd18, 3'b111};	// Note: 4A#Bb
	assign memory[	 60	] =	{1'b0, 6'd29, 6'd18, 3'b111};	// Note: 3C#Db
	assign memory[	 61	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	 62	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	 63	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	 64	] =	{1'b0, 6'd29, 6'd6, 3'b111};	// Note: 3C#Db
	assign memory[	 65	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 66	] =	{1'b0, 6'd38, 6'd36, 3'b111};	// Note: 4A#Bb
	assign memory[	 67	] =	{1'b0, 6'd29, 6'd36, 3'b111};	// Note: 3C#Db
	assign memory[	 68	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 69	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 70	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 71	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 72	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 73	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 74	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	 75	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	 76	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	 77	] =	{1'b0, 6'd29, 6'd6, 3'b111};	// Note: 3C#Db
	assign memory[	 78	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 79	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	 80	] =	{1'b0, 6'd29, 6'd6, 3'b111};	// Note: 3C#Db
	assign memory[	 81	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	 82	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 83	] =	{1'b0, 6'd29, 6'd8, 3'b111};	// Note: 3C#Db
	assign memory[	 84	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 85	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 86	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 87	] =	{1'b0, 6'd29, 6'd8, 3'b111};	// Note: 3C#Db
	assign memory[	 88	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 89	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 90	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	 91	] =	{1'b0, 6'd29, 6'd8, 3'b111};	// Note: 3C#Db
	assign memory[	 92	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	 93	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	 94	] =	{1'b0, 6'd38, 6'd12, 3'b111};	// Note: 4A#Bb
	assign memory[	 95	] =	{1'b0, 6'd29, 6'd12, 3'b111};	// Note: 3C#Db
	assign memory[	 96	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	 97	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	 98	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	 99	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	100	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	101	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	102	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	103	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	104	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	105	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	106	] =	{1'b0, 6'd9, 6'd24, 3'b111};	// Note: 1F
	assign memory[	107	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	108	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	109	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	110	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	111	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	112	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	113	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	114	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	115	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	116	] =	{1'b0, 6'd9, 6'd24, 3'b111};	// Note: 1F
	assign memory[	117	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	118	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	119	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	120	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	121	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	122	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	123	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	124	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	125	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	126	] =	{1'b0, 6'd11, 6'd12, 3'b111};	// Note: 1G
	assign memory[	127	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	128	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	129	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	130	] =	{1'b0, 6'd13, 6'd12, 3'b111};	// Note: 2A
	assign memory[	131	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	132	] =	{1'b0, 6'd38, 6'd24, 3'b111};	// Note: 4A#Bb
	assign memory[	133	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	134	] =	{1'b0, 6'd14, 6'd24, 3'b111};	// Note: 2A#Bb
	assign memory[	135	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	136	] =	{1'b0, 6'd33, 6'd36, 3'b111};	// Note: 3F
	assign memory[	137	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	138	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Db
	assign memory[	139	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	140	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	141	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Db
	assign memory[	142	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	143	] =	{1'b0, 6'd28, 6'd8, 3'b111};	// Note: 3C
	assign memory[	144	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	145	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	146	] =	{1'b0, 6'd30, 6'd18, 3'b111};	// Note: 3D
	assign memory[	147	] =	{1'b0, 6'd14, 6'd24, 3'b111};	// Note: 2A#Bb
	assign memory[	148	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	149	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	150	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	151	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	152	] =	{1'b0, 6'd30, 6'd6, 3'b111};	// Note: 3D
	assign memory[	153	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	154	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	155	] =	{1'b0, 6'd30, 6'd6, 3'b111};	// Note: 3D
	assign memory[	156	] =	{1'b0, 6'd14, 6'd24, 3'b111};	// Note: 2A#Bb
	assign memory[	157	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	158	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	159	] =	{1'b0, 6'd31, 6'd6, 3'b111};	// Note: 3D#Eb
	assign memory[	160	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	161	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	162	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	163	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	164	] =	{1'b0, 6'd43, 6'd6, 3'b111};	// Note: 4D#Eb
	assign memory[	165	] =	{1'b0, 6'd35, 6'd6, 3'b111};	// Note: 3G
	assign memory[	166	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	167	] =	{1'b0, 6'd45, 6'd48, 3'b111};	// Note: 4F
	assign memory[	168	] =	{1'b0, 6'd36, 6'd18, 3'b111};	// Note: 3G#Ab
	assign memory[	169	] =	{1'b0, 6'd12, 6'd24, 3'b111};	// Note: 1G#Ab
	assign memory[	170	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	171	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	172	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	173	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	174	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	175	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	176	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	177	] =	{1'b1, 6'd0, 6'd2, 3'b111};	// Note: rest
	assign memory[	178	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	179	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	180	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	181	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	182	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	183	] =	{1'b1, 6'd0, 6'd2, 3'b111};	// Note: rest
	assign memory[	184	] =	{1'b0, 6'd43, 6'd6, 3'b111};	// Note: 4D#Eb
	assign memory[	185	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	186	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	187	] =	{1'b0, 6'd12, 6'd24, 3'b111};	// Note: 1G#Ab
	assign memory[	188	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	189	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	190	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	191	] =	{1'b0, 6'd45, 6'd8, 3'b111};	// Note: 4F
	assign memory[	192	] =	{1'b0, 6'd36, 6'd8, 3'b111};	// Note: 3G#Ab
	assign memory[	193	] =	{1'b0, 6'd12, 6'd24, 3'b111};	// Note: 1G#Ab
	assign memory[	194	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	195	] =	{1'b0, 6'd46, 6'd8, 3'b111};	// Note: 4F#Gb
	assign memory[	196	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	197	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	198	] =	{1'b0, 6'd48, 6'd8, 3'b111};	// Note: 4G#Ab
	assign memory[	199	] =	{1'b0, 6'd40, 6'd8, 3'b111};	// Note: 4C
	assign memory[	200	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	201	] =	{1'b0, 6'd50, 6'd48, 3'b111};	// Note: 5A#Bb
	assign memory[	202	] =	{1'b0, 6'd41, 6'd36, 3'b111};	// Note: 4C#Db
	assign memory[	203	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	204	] =	{1'b1, 6'd0, 6'd36, 3'b111};	// Note: rest
	assign memory[	205	] =	{1'b0, 6'd34, 6'd6, 3'b111};	// Note: 3F#Gb
	assign memory[	206	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	207	] =	{1'b0, 6'd34, 6'd6, 3'b111};	// Note: 3F#Gb
	assign memory[	208	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	209	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	210	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	211	] =	{1'b1, 6'd0, 6'd2, 3'b111};	// Note: rest
	assign memory[	212	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	213	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	214	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	215	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	216	] =	{1'b0, 6'd8, 6'd8, 3'b111};	// Note: 1E
	assign memory[	217	] =	{1'b1, 6'd0, 6'd2, 3'b111};	// Note: rest
	assign memory[	218	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	219	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	220	] =	{1'b0, 6'd50, 6'd9, 3'b111};	// Note: 5A#Bb
	assign memory[	221	] =	{1'b0, 6'd41, 6'd12, 3'b111};	// Note: 4C#Db
	assign memory[	222	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	223	] =	{1'b1, 6'd0, 6'd9, 3'b111};	// Note: rest
	assign memory[	224	] =	{1'b0, 6'd50, 6'd9, 3'b111};	// Note: 5A#Bb
	assign memory[	225	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	226	] =	{1'b0, 6'd41, 6'd12, 3'b111};	// Note: 4C#Db
	assign memory[	227	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	228	] =	{1'b0, 6'd50, 6'd6, 3'b111};	// Note: 5A#Bb
	assign memory[	229	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	230	] =	{1'b0, 6'd50, 6'd8, 3'b111};	// Note: 5A#Bb
	assign memory[	231	] =	{1'b0, 6'd41, 6'd8, 3'b111};	// Note: 4C#Db
	assign memory[	232	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	233	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	234	] =	{1'b0, 6'd48, 6'd8, 3'b111};	// Note: 4G#Ab
	assign memory[	235	] =	{1'b0, 6'd40, 6'd8, 3'b111};	// Note: 4C
	assign memory[	236	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	237	] =	{1'b0, 6'd46, 6'd8, 3'b111};	// Note: 4F#Gb
	assign memory[	238	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	239	] =	{1'b0, 6'd17, 6'd8, 3'b111};	// Note: rest
	assign memory[	240	] =	{1'b0, 6'd41, 6'd24, 3'b111};	// Note: 2C#Db
	assign memory[	241	] =	{1'b0, 6'd48, 6'd18, 3'b111};	// Note: 4C#Db
	assign memory[	242	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: 4G#Ab
	assign memory[	243	] =	{1'b0, 6'd46, 6'd18, 3'b111};	// Note: rest
	assign memory[	244	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 4F#Gb
	assign memory[	245	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	246	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: rest
	assign memory[	247	] =	{1'b0, 6'd36, 6'd48, 3'b111};	// Note: 4F
	assign memory[	248	] =	{1'b0, 6'd17, 6'd8, 3'b111};	// Note: 3G#Ab
	assign memory[	249	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: 2C#Db
	assign memory[	250	] =	{1'b0, 6'd36, 6'd8, 3'b111};	// Note: rest
	assign memory[	251	] =	{1'b0, 6'd17, 6'd8, 3'b111};	// Note: 3G#Ab
	assign memory[	252	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: 2C#Db
	assign memory[	253	] =	{1'b0, 6'd34, 6'd8, 3'b111};	// Note: rest
	assign memory[	254	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 3F#Gb
	assign memory[	255	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: 2B
	assign memory[	256	] =	{1'b0, 6'd17, 6'd24, 3'b111};	// Note: 2C#Db
	assign memory[	257	] =	{1'b0, 6'd36, 6'd18, 3'b111};	// Note: 3G#Ab
	assign memory[	258	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	259	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	260	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	261	] =	{1'b0, 6'd45, 6'd24, 3'b111};	// Note: 4F
	assign memory[	262	] =	{1'b0, 6'd17, 6'd24, 3'b111};	// Note: 2C#Db
	assign memory[	263	] =	{1'b0, 6'd36, 6'd24, 3'b111};	// Note: 3G#Ab
	assign memory[	264	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	265	] =	{1'b0, 6'd34, 6'd8, 3'b111};	// Note: 3F#Gb
	assign memory[	266	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	267	] =	{1'b0, 6'd36, 6'd8, 3'b111};	// Note: 3G#Ab
	assign memory[	268	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	269	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	270	] =	{1'b0, 6'd34, 6'd24, 3'b111};	// Note: 3F#Gb
	assign memory[	271	] =	{1'b0, 6'd43, 6'd12, 3'b111};	// Note: 4D#Eb
	assign memory[	272	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	273	] =	{1'b0, 6'd43, 6'd12, 3'b111};	// Note: 4D#Eb
	assign memory[	274	] =	{1'b0, 6'd34, 6'd6, 3'b111};	// Note: 3F#Gb
	assign memory[	275	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	276	] =	{1'b0, 6'd34, 6'd4, 3'b111};	// Note: 3F#Gb
	assign memory[	277	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	278	] =	{1'b0, 6'd45, 6'd2, 3'b111};	// Note: 4F
	assign memory[	279	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	280	] =	{1'b0, 6'd33, 6'd2, 3'b111};	// Note: 3F
	assign memory[	281	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	282	] =	{1'b0, 6'd46, 6'd4, 3'b111};	// Note: 4F#Gb
	assign memory[	283	] =	{1'b0, 6'd34, 6'd48, 3'b111};	// Note: 3F#Gb
	assign memory[	284	] =	{1'b0, 6'd15, 6'd12, 3'b111};	// Note: 2B
	assign memory[	285	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	286	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	287	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	288	] =	{1'b0, 6'd34, 6'd4, 3'b111};	// Note: 3F#Gb
	assign memory[	289	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	290	] =	{1'b0, 6'd14, 6'd4, 3'b111};	// Note: 2A#Bb
	assign memory[	291	] =	{1'b0, 6'd34, 6'd8, 3'b111};	// Note: 3F#Gb
	assign memory[	292	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	293	] =	{1'b0, 6'd36, 6'd4, 3'b111};	// Note: 3G#Ab
	assign memory[	294	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	295	] =	{1'b0, 6'd38, 6'd4, 3'b111};	// Note: 4A#Bb
	assign memory[	296	] =	{1'b0, 6'd15, 6'd24, 3'b111};	// Note: 2B
	assign memory[	297	] =	{1'b0, 6'd36, 6'd24, 3'b111};	// Note: 3G#Ab
	assign memory[	298	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	299	] =	{1'b0, 6'd15, 6'd12, 3'b111};	// Note: 2B
	assign memory[	300	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	301	] =	{1'b0, 6'd15, 6'd8, 3'b111};	// Note: 2B
	assign memory[	302	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	303	] =	{1'b0, 6'd34, 6'd4, 3'b111};	// Note: 3F#Gb
	assign memory[	304	] =	{1'b0, 6'd43, 6'd12, 3'b111};	// Note: 4D#Eb
	assign memory[	305	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	306	] =	{1'b0, 6'd15, 6'd4, 3'b111};	// Note: 2B
	assign memory[	307	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	308	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	309	] =	{1'b0, 6'd33, 6'd24, 3'b111};	// Note: 3F
	assign memory[	310	] =	{1'b0, 6'd41, 6'd12, 3'b111};	// Note: 4C#Db
	assign memory[	311	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	312	] =	{1'b0, 6'd41, 6'd12, 3'b111};	// Note: 4C#Db
	assign memory[	313	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	314	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	315	] =	{1'b0, 6'd33, 6'd4, 3'b111};	// Note: 3F
	assign memory[	316	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	317	] =	{1'b0, 6'd43, 6'd2, 3'b111};	// Note: 4D#Eb
	assign memory[	318	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	319	] =	{1'b0, 6'd31, 6'd2, 3'b111};	// Note: 3D#Eb
	assign memory[	320	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	321	] =	{1'b0, 6'd45, 6'd4, 3'b111};	// Note: 4F
	assign memory[	322	] =	{1'b0, 6'd33, 6'd48, 3'b111};	// Note: 3F
	assign memory[	323	] =	{1'b0, 6'd14, 6'd12, 3'b111};	// Note: 2A#Bb
	assign memory[	324	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	325	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	326	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	327	] =	{1'b0, 6'd21, 6'd4, 3'b111};	// Note: 2F
	assign memory[	328	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	329	] =	{1'b0, 6'd21, 6'd4, 3'b111};	// Note: 2F
	assign memory[	330	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	331	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	332	] =	{1'b0, 6'd34, 6'd4, 3'b111};	// Note: 3F#Gb
	assign memory[	333	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	334	] =	{1'b0, 6'd14, 6'd4, 3'b111};	// Note: 2A#Bb
	assign memory[	335	] =	{1'b0, 6'd36, 6'd24, 3'b111};	// Note: 3G#Ab
	assign memory[	336	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	337	] =	{1'b0, 6'd35, 6'd24, 3'b111};	// Note: 3G
	assign memory[	338	] =	{1'b0, 6'd43, 6'd12, 3'b111};	// Note: 4D#Eb
	assign memory[	339	] =	{1'b0, 6'd14, 6'd12, 3'b111};	// Note: 2A#Bb
	assign memory[	340	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	341	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	342	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	343	] =	{1'b0, 6'd33, 6'd4, 3'b111};	// Note: 3F
	assign memory[	344	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	345	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	346	] =	{1'b0, 6'd14, 6'd4, 3'b111};	// Note: 2A#Bb
	assign memory[	347	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	348	] =	{1'b0, 6'd16, 6'd8, 3'b111};	// Note: 2C
	assign memory[	349	] =	{1'b0, 6'd32, 6'd24, 3'b111};	// Note: 3E
	assign memory[	350	] =	{1'b0, 6'd40, 6'd24, 3'b111};	// Note: 4C
	assign memory[	351	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	352	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	353	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	354	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	355	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	356	] =	{1'b0, 6'd44, 6'd6, 3'b111};	// Note: 4E
	assign memory[	357	] =	{1'b0, 6'd32, 6'd48, 3'b111};	// Note: 3E
	assign memory[	358	] =	{1'b0, 6'd16, 6'd18, 3'b111};	// Note: 2C
	assign memory[	359	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	360	] =	{1'b0, 6'd16, 6'd8, 3'b111};	// Note: 2C
	assign memory[	361	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	362	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	363	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	364	] =	{1'b0, 6'd33, 6'd4, 3'b111};	// Note: 3F
	assign memory[	365	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	366	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	367	] =	{1'b0, 6'd35, 6'd24, 3'b111};	// Note: 3G
	assign memory[	368	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	369	] =	{1'b0, 6'd35, 6'd12, 3'b111};	// Note: 3G
	assign memory[	370	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	371	] =	{1'b0, 6'd35, 6'd4, 3'b111};	// Note: 3G
	assign memory[	372	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	373	] =	{1'b0, 6'd37, 6'd4, 3'b111};	// Note: 4A
	assign memory[	374	] =	{1'b1, 6'd0, 6'd4, 3'b111};	// Note: rest
	assign memory[	375	] =	{1'b0, 6'd47, 6'd4, 3'b111};	// Note: 4G
	assign memory[	376	] =	{1'b0, 6'd38, 6'd24, 3'b111};	// Note: 4A#Bb
	assign memory[	377	] =	{1'b0, 6'd16, 6'd12, 3'b111};	// Note: 2C
	assign memory[	378	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	379	] =	{1'b0, 6'd16, 6'd8, 3'b111};	// Note: 2C
	assign memory[	380	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	381	] =	{1'b0, 6'd40, 6'd4, 3'b111};	// Note: 4C
	assign memory[	382	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	383	] =	{1'b0, 6'd16, 6'd4, 3'b111};	// Note: 2C
	assign memory[	384	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	385	] =	{1'b0, 6'd9, 6'd8, 3'b111};	// Note: 1F
	assign memory[	386	] =	{1'b0, 6'd37, 6'd24, 3'b111};	// Note: 4A
	assign memory[	387	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	388	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	389	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	390	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	391	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	392	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	393	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	394	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	395	] =	{1'b0, 6'd9, 6'd6, 3'b111};	// Note: 1F
	assign memory[	396	] =	{1'b0, 6'd33, 6'd24, 3'b111};	// Note: 3F
	assign memory[	397	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	398	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	399	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	400	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	401	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	402	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	403	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	404	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	405	] =	{1'b0, 6'd9, 6'd6, 3'b111};	// Note: 1F
	assign memory[	406	] =	{1'b0, 6'd33, 6'd24, 3'b111};	// Note: 3F
	assign memory[	407	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	408	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	409	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	410	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	411	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	412	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	413	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	414	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	415	] =	{1'b0, 6'd11, 6'd6, 3'b111};	// Note: 1G
	assign memory[	416	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	417	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	418	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	419	] =	{1'b0, 6'd13, 6'd12, 3'b111};	// Note: 2A
	assign memory[	420	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	421	] =	{1'b0, 6'd25, 6'd12, 3'b111};	// Note: 3A
	assign memory[	422	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	423	] =	{1'b0, 6'd14, 6'd12, 3'b111};	// Note: 2A#Bb
	assign memory[	424	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	425	] =	{1'b0, 6'd38, 6'd24, 3'b111};	// Note: 4A#Bb
	assign memory[	426	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	427	] =	{1'b0, 6'd33, 6'd24, 3'b111};	// Note: 3F
	assign memory[	428	] =	{1'b0, 6'd14, 6'd36, 3'b111};	// Note: 2A#Bb
	assign memory[	429	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	430	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	431	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	432	] =	{1'b0, 6'd30, 6'd8, 3'b111};	// Note: 3D
	assign memory[	433	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	434	] =	{1'b0, 6'd12, 6'd8, 3'b111};	// Note: 1G#Ab
	assign memory[	435	] =	{1'b0, 6'd28, 6'd8, 3'b111};	// Note: 3C
	assign memory[	436	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	437	] =	{1'b0, 6'd14, 6'd8, 3'b111};	// Note: 2A#Bb
	assign memory[	438	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	439	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	440	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	441	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	442	] =	{1'b0, 6'd30, 6'd6, 3'b111};	// Note: 3D
	assign memory[	443	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	444	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	445	] =	{1'b0, 6'd14, 6'd6, 3'b111};	// Note: 2A#Bb
	assign memory[	446	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	447	] =	{1'b0, 6'd38, 6'd6, 3'b111};	// Note: 4A#Bb
	assign memory[	448	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	449	] =	{1'b0, 6'd31, 6'd6, 3'b111};	// Note: 3D#Eb
	assign memory[	450	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	451	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	452	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	453	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	454	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	455	] =	{1'b0, 6'd35, 6'd6, 3'b111};	// Note: 3G
	assign memory[	456	] =	{1'b0, 6'd43, 6'd6, 3'b111};	// Note: 4D#Eb
	assign memory[	457	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	458	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: 4F
	assign memory[	459	] =	{1'b0, 6'd12, 6'd48, 3'b111};	// Note: 1G#Ab
	assign memory[	460	] =	{1'b0, 6'd36, 6'd24, 3'b111};	// Note: 3G#Ab
	assign memory[	461	] =	{1'b1, 6'd0, 6'd18, 3'b111};	// Note: rest
	assign memory[	462	] =	{1'b0, 6'd38, 6'd18, 3'b111};	// Note: 4A#Bb
	assign memory[	463	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	464	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	465	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	466	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	467	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	468	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	469	] =	{1'b0, 6'd12, 6'd2, 3'b111};	// Note: 1G#Ab
	assign memory[	470	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	471	] =	{1'b0, 6'd42, 6'd4, 3'b111};	// Note: 4D
	assign memory[	472	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	473	] =	{1'b0, 6'd10, 6'd4, 3'b111};	// Note: 1F#Gb
	assign memory[	474	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	475	] =	{1'b0, 6'd43, 6'd2, 3'b111};	// Note: 4D#Eb
	assign memory[	476	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	477	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	478	] =	{1'b0, 6'd45, 6'd24, 3'b111};	// Note: 4F
	assign memory[	479	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	480	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	481	] =	{1'b0, 6'd45, 6'd12, 3'b111};	// Note: 4F
	assign memory[	482	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	483	] =	{1'b0, 6'd12, 6'd12, 3'b111};	// Note: 1G#Ab
	assign memory[	484	] =	{1'b0, 6'd36, 6'd24, 3'b111};	// Note: 3G#Ab
	assign memory[	485	] =	{1'b0, 6'd45, 6'd8, 3'b111};	// Note: 4F
	assign memory[	486	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	487	] =	{1'b0, 6'd38, 6'd8, 3'b111};	// Note: 4A#Bb
	assign memory[	488	] =	{1'b0, 6'd46, 6'd8, 3'b111};	// Note: 4F#Gb
	assign memory[	489	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	490	] =	{1'b0, 6'd40, 6'd8, 3'b111};	// Note: 4C
	assign memory[	491	] =	{1'b0, 6'd48, 6'd8, 3'b111};	// Note: 4G#Ab
	assign memory[	492	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	493	] =	{1'b0, 6'd41, 6'd8, 3'b111};	// Note: 4C#Db
	assign memory[	494	] =	{1'b0, 6'd50, 6'd24, 3'b111};	// Note: 5A#Bb
	assign memory[	495	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	496	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	497	] =	{1'b0, 6'd41, 6'd24, 3'b111};	// Note: 4C#Db
	assign memory[	498	] =	{1'b0, 6'd50, 6'd48, 3'b111};	// Note: 5A#Bb
	assign memory[	499	] =	{1'b0, 6'd10, 6'd48, 3'b111};	// Note: 1F#Gb
	assign memory[	500	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	501	] =	{1'b0, 6'd8, 6'd8, 3'b111};	// Note: 1E
	assign memory[	502	] =	{1'b1, 6'd0, 6'd8, 3'b111};	// Note: rest
	assign memory[	503	] =	{1'b0, 6'd10, 6'd8, 3'b111};	// Note: 1F#Gb
	assign memory[	504	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	505	] =	{1'b0, 6'd10, 6'd24, 3'b111};	// Note: 1F#Gb
	assign memory[	506	] =	{1'b0, 6'd44, 6'd24, 3'b111};	// Note: 4E
	assign memory[	507	] =	{1'b0, 6'd53, 6'd24, 3'b111};	// Note: 5C#Db
	assign memory[	508	] =	{1'b1, 6'd0, 6'd22, 3'b111};	// Note: rest
	assign memory[	509	] =	{1'b0, 6'd44, 6'd24, 3'b111};	// Note: 4E
	assign memory[	510	] =	{1'b0, 6'd53, 6'd24, 3'b111};	// Note: 5C#Db
	assign memory[	511	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest

	SONG 2

	assign memory[	512	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	513	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	514	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	515	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	516	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	517	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: res
	assign memory[	518	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	519	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	520	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	521	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	522	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	523	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	524	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	525	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	526	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	527	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	528	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	529	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	530	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	531	] =	{1'b0, 6'd44, 6'd3, 3'b111};	// Note: 4E
	assign memory[	532	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	533	] =	{1'b0, 6'd42, 6'd3, 3'b111};	// Note: 4D
	assign memory[	534	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	535	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	536	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	537	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	538	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	539	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	540	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	541	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	542	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	543	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	544	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	545	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	546	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	547	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	548	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	549	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	550	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	551	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	552	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	553	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	554	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	555	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	556	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	557	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	558	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	559	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	560	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	561	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	562	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	563	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	564	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	565	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	566	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	567	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	568	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	569	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	570	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	571	] =	{1'b0, 6'd39, 6'd18, 3'b111};	// Note: 4B
	assign memory[	572	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	573	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	574	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	575	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	576	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	577	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	578	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	579	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	580	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	581	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	582	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	583	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	584	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	585	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	586	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	587	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	588	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	589	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	590	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	591	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	592	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	593	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	594	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	595	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	596	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	597	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	598	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	599	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	600	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	601	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	602	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	603	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	604	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	605	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	606	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	607	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	608	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	609	] =	{1'b0, 6'd32, 6'd24, 3'b111};	// Note: 3E
	assign memory[	610	] =	{1'b0, 6'd37, 6'd24, 3'b111};	// Note: 4A
	assign memory[	611	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	612	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	613	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	614	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	615	] =	{1'b0, 6'd15, 6'd6, 3'b111};	// Note: 2B
	assign memory[	616	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	617	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	618	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	619	] =	{1'b0, 6'd18, 6'd6, 3'b111};	// Note: 2D
	assign memory[	620	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	621	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	622	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	623	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	624	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	625	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	626	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	627	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: 4F
	assign memory[	628	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	629	] =	{1'b0, 6'd49, 6'd12, 3'b111};	// Note: 5A
	assign memory[	630	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	631	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	632	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	633	] =	{1'b0, 6'd40, 6'd3, 3'b111};	// Note: 4C
	assign memory[	634	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	635	] =	{1'b0, 6'd40, 6'd3, 3'b111};	// Note: 4C
	assign memory[	636	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	637	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	638	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	639	] =	{1'b0, 6'd47, 6'd6, 3'b111};	// Note: 4G
	assign memory[	640	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	641	] =	{1'b0, 6'd9, 6'd6, 3'b111};	// Note: 1F
	assign memory[	642	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	643	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: 4F
	assign memory[	644	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	645	] =	{1'b0, 6'd35, 6'd18, 3'b111};	// Note: 3G
	assign memory[	646	] =	{1'b0, 6'd44, 6'd18, 3'b111};	// Note: 4E
	assign memory[	647	] =	{1'b0, 6'd4, 6'd6, 3'b111};	// Note: 1C
	assign memory[	648	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	649	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	650	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	651	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	652	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	653	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	654	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	655	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	656	] =	{1'b0, 6'd4, 6'd6, 3'b111};	// Note: 1C
	assign memory[	657	] =	{1'b0, 6'd35, 6'd6, 3'b111};	// Note: 3G
	assign memory[	658	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	659	] =	{1'b0, 6'd11, 6'd6, 3'b111};	// Note: 1G
	assign memory[	660	] =	{1'b0, 6'd37, 6'd3, 3'b111};	// Note: 4A
	assign memory[	661	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	662	] =	{1'b0, 6'd35, 6'd3, 3'b111};	// Note: 3G
	assign memory[	663	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	664	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	665	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	666	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	667	] =	{1'b0, 6'd11, 6'd6, 3'b111};	// Note: 1G
	assign memory[	668	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	669	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	670	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	671	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	672	] =	{1'b0, 6'd15, 6'd6, 3'b111};	// Note: 2B
	assign memory[	673	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	674	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	675	] =	{1'b0, 6'd27, 6'd6, 3'b111};	// Note: 3B
	assign memory[	676	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	677	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	678	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	679	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	680	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	681	] =	{1'b0, 6'd27, 6'd6, 3'b111};	// Note: 3B
	assign memory[	682	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	683	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	684	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	685	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	686	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	687	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	688	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	689	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	690	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	691	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	692	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	693	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	694	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	695	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	696	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	697	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	698	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	699	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	700	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	701	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	702	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	703	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	704	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	705	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	706	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	707	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	708	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	709	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	710	] =	{1'b0, 6'd13, 6'd12, 3'b111};	// Note: 2A
	assign memory[	711	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	712	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	713	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	714	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	715	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	716	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	717	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	718	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	719	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	720	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	721	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	722	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	723	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	724	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	725	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	726	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	727	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	728	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	729	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	730	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	731	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	732	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	733	] =	{1'b0, 6'd44, 6'd3, 3'b111};	// Note: 4E
	assign memory[	734	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	735	] =	{1'b0, 6'd42, 6'd3, 3'b111};	// Note: 4D
	assign memory[	736	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	737	] =	{1'b0, 6'd8, 6'd6, 3'b111};	// Note: 1E
	assign memory[	738	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	739	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	740	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	741	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	742	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	743	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	744	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	745	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	746	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	747	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	748	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	749	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	750	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	751	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	752	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	753	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	754	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	755	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	756	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	757	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	758	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	759	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	760	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	761	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	762	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	763	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	764	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	765	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	766	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	767	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	768	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	769	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	770	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	771	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	772	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	773	] =	{1'b0, 6'd39, 6'd18, 3'b111};	// Note: 4B
	assign memory[	774	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	775	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	776	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	777	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	778	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	779	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	780	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	781	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	782	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	783	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	784	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	785	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	786	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	787	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	788	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	789	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	790	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	791	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	792	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	793	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	794	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	795	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	796	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	797	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	798	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	799	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	800	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	801	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	802	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	803	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	804	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	805	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	806	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	807	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	808	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	809	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	810	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	811	] =	{1'b0, 6'd32, 6'd24, 3'b111};	// Note: 3E
	assign memory[	812	] =	{1'b0, 6'd37, 6'd24, 3'b111};	// Note: 4A
	assign memory[	813	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	814	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	815	] =	{1'b0, 6'd25, 6'd6, 3'b111};	// Note: 3A
	assign memory[	816	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	817	] =	{1'b0, 6'd15, 6'd6, 3'b111};	// Note: 2B
	assign memory[	818	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	819	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	820	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	821	] =	{1'b0, 6'd18, 6'd6, 3'b111};	// Note: 2D
	assign memory[	822	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	823	] =	{1'b0, 6'd33, 6'd12, 3'b111};	// Note: 3F
	assign memory[	824	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	825	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	826	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	827	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	828	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	829	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: 4F
	assign memory[	830	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	831	] =	{1'b0, 6'd49, 6'd12, 3'b111};	// Note: 5A
	assign memory[	832	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	833	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	834	] =	{1'b0, 6'd6, 6'd6, 3'b111};	// Note: 1D
	assign memory[	835	] =	{1'b0, 6'd40, 6'd3, 3'b111};	// Note: 4C
	assign memory[	836	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	837	] =	{1'b0, 6'd40, 6'd3, 3'b111};	// Note: 4C
	assign memory[	838	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	839	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	840	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	841	] =	{1'b0, 6'd47, 6'd6, 3'b111};	// Note: 4G
	assign memory[	842	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	843	] =	{1'b0, 6'd9, 6'd6, 3'b111};	// Note: 1F
	assign memory[	844	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	845	] =	{1'b0, 6'd45, 6'd6, 3'b111};	// Note: 4F
	assign memory[	846	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	847	] =	{1'b0, 6'd35, 6'd18, 3'b111};	// Note: 3G
	assign memory[	848	] =	{1'b0, 6'd44, 6'd18, 3'b111};	// Note: 4E
	assign memory[	849	] =	{1'b0, 6'd4, 6'd6, 3'b111};	// Note: 1C
	assign memory[	850	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	851	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	852	] =	{1'b1, 6'd0, 6'd12, 3'b111};	// Note: rest
	assign memory[	853	] =	{1'b0, 6'd16, 6'd6, 3'b111};	// Note: 2C
	assign memory[	854	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	855	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	856	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	857	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	858	] =	{1'b0, 6'd4, 6'd6, 3'b111};	// Note: 1C
	assign memory[	859	] =	{1'b0, 6'd35, 6'd6, 3'b111};	// Note: 3G
	assign memory[	860	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	861	] =	{1'b0, 6'd11, 6'd6, 3'b111};	// Note: 1G
	assign memory[	862	] =	{1'b0, 6'd37, 6'd3, 3'b111};	// Note: 4A
	assign memory[	863	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	864	] =	{1'b0, 6'd35, 6'd3, 3'b111};	// Note: 3G
	assign memory[	865	] =	{1'b1, 6'd0, 6'd3, 3'b111};	// Note: rest
	assign memory[	866	] =	{1'b0, 6'd33, 6'd6, 3'b111};	// Note: 3F
	assign memory[	867	] =	{1'b0, 6'd42, 6'd6, 3'b111};	// Note: 4D
	assign memory[	868	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	869	] =	{1'b0, 6'd11, 6'd6, 3'b111};	// Note: 1G
	assign memory[	870	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	871	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	872	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	873	] =	{1'b0, 6'd39, 6'd12, 3'b111};	// Note: 4B
	assign memory[	874	] =	{1'b0, 6'd15, 6'd6, 3'b111};	// Note: 2B
	assign memory[	875	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	876	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	877	] =	{1'b0, 6'd27, 6'd6, 3'b111};	// Note: 3B
	assign memory[	878	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	879	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	880	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	881	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	882	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	883	] =	{1'b0, 6'd27, 6'd6, 3'b111};	// Note: 3B
	assign memory[	884	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	885	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	886	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	887	] =	{1'b0, 6'd42, 6'd12, 3'b111};	// Note: 4D
	assign memory[	888	] =	{1'b0, 6'd39, 6'd6, 3'b111};	// Note: 4B
	assign memory[	889	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	890	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	891	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	892	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	893	] =	{1'b0, 6'd44, 6'd12, 3'b111};	// Note: 4E
	assign memory[	894	] =	{1'b0, 6'd40, 6'd6, 3'b111};	// Note: 4C
	assign memory[	895	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	896	] =	{1'b0, 6'd24, 6'd6, 3'b111};	// Note: 2G#Ab
	assign memory[	897	] =	{1'b0, 6'd36, 6'd6, 3'b111};	// Note: 3G#Ab
	assign memory[	898	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	899	] =	{1'b0, 6'd40, 6'd12, 3'b111};	// Note: 4C
	assign memory[	900	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	901	] =	{1'b0, 6'd37, 6'd6, 3'b111};	// Note: 4A
	assign memory[	902	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	903	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	904	] =	{1'b0, 6'd32, 6'd6, 3'b111};	// Note: 3E
	assign memory[	905	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	906	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	907	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	908	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	909	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	910	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	911	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	912	] =	{1'b0, 6'd13, 6'd12, 3'b111};	// Note: 2A
	assign memory[	913	] =	{1'b0, 6'd32, 6'd12, 3'b111};	// Note: 3E
	assign memory[	914	] =	{1'b0, 6'd37, 6'd12, 3'b111};	// Note: 4A
	assign memory[	915	] =	{1'b1, 6'd0, 6'd24, 3'b111};	// Note: rest
	assign memory[	916	] =	{1'b0, 6'd28, 6'd24, 3'b111};	// Note: 3C
	assign memory[	917	] =	{1'b0, 6'd32, 6'd24, 3'b111};	// Note: 3E
	assign memory[	918	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	919	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	920	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	921	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	922	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	923	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	924	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	925	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	926	] =	{1'b0, 6'd25, 6'd24, 3'b111};	// Note: 3A
	assign memory[	927	] =	{1'b0, 6'd28, 6'd24, 3'b111};	// Note: 3C
	assign memory[	928	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	929	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	930	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	931	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	932	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	933	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	934	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	935	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	936	] =	{1'b0, 6'd27, 6'd24, 3'b111};	// Note: 3B
	assign memory[	937	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	938	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	939	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	940	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	941	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	942	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	943	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	944	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	945	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	946	] =	{1'b0, 6'd24, 6'd24, 3'b111};	// Note: 2G#Ab
	assign memory[	947	] =	{1'b0, 6'd27, 6'd24, 3'b111};	// Note: 3B
	assign memory[	948	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	949	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	950	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	951	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	952	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	953	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	954	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	955	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	956	] =	{1'b0, 6'd25, 6'd24, 3'b111};	// Note: 3A
	assign memory[	957	] =	{1'b0, 6'd28, 6'd24, 3'b111};	// Note: 3C
	assign memory[	958	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	959	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	960	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	961	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	962	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	963	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	964	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	965	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	966	] =	{1'b0, 6'd20, 6'd24, 3'b111};	// Note: 2E
	assign memory[	967	] =	{1'b0, 6'd25, 6'd24, 3'b111};	// Note: 3A
	assign memory[	968	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	969	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	970	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	971	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	972	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	973	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	974	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	975	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	976	] =	{1'b0, 6'd24, 6'd24, 3'b111};	// Note: 2G#Ab
	assign memory[	977	] =	{1'b0, 6'd20, 6'd24, 3'b111};	// Note: 2E
	assign memory[	978	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	979	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	980	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	981	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	982	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	983	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	984	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	985	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	986	] =	{1'b0, 6'd24, 6'd24, 3'b111};	// Note: 2G#Ab
	assign memory[	987	] =	{1'b0, 6'd27, 6'd24, 3'b111};	// Note: 3B
	assign memory[	988	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	989	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	990	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	991	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	992	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	993	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	994	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	995	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	996	] =	{1'b0, 6'd28, 6'd24, 3'b111};	// Note: 3C
	assign memory[	997	] =	{1'b0, 6'd32, 6'd24, 3'b111};	// Note: 3E
	assign memory[	998	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	999	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1000	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	1001	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1002	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	1003	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1004	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	1005	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1006	] =	{1'b0, 6'd25, 6'd24, 3'b111};	// Note: 3A
	assign memory[	1007	] =	{1'b0, 6'd28, 6'd24, 3'b111};	// Note: 3C
	assign memory[	1008	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	1009	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1010	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	1011	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1012	] =	{1'b0, 6'd13, 6'd6, 3'b111};	// Note: 2A
	assign memory[	1013	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1014	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	1015	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1016	] =	{1'b0, 6'd30, 6'd24, 3'b111};	// Note: 3D
	assign memory[	1017	] =	{1'b0, 6'd27, 6'd24, 3'b111};	// Note: 3B
	assign memory[	1018	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	1019	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1020	] =	{1'b0, 6'd20, 6'd6, 3'b111};	// Note: 2E
	assign memory[	1021	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest
	assign memory[	1022	] =	{1'b0, 6'd12, 6'd6, 3'b111};	// Note: 1G#Ab
	assign memory[	1023	] =	{1'b1, 6'd0, 6'd6, 3'b111};	// Note: rest

// Song 3

	assign memory[	1024	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1025	] =	{1'b0, 6'd24, 6'd18, 3'd4};	// Note: 2G#Ab
	assign memory[	1026	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1027	] =	{1'b0, 6'd39, 6'd3, 3'd3};	// Note: 4B
	assign memory[	1028	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1029	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1030	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1031	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1032	] =	{1'b0, 6'd24, 6'd6, 3'd4};	// Note: 2G#Ab
	assign memory[	1033	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1034	] =	{1'b0, 6'd24, 6'd18, 3'd4};	// Note: 2G#Ab
	assign memory[	1035	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1036	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1037	] =	{1'b0, 6'd31, 6'd3, 3'd3};	// Note: 3D#Eb
	assign memory[	1038	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1039	] =	{1'b0, 6'd31, 6'd6, 3'd5};	// Note: 3D#Eb
	assign memory[	1040	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1041	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1042	] =	{1'b0, 6'd24, 6'd6, 3'd4};	// Note: 2G#Ab
	assign memory[	1043	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1044	] =	{1'b0, 6'd22, 6'd24, 3'd4};	// Note: 2F#Gb
	assign memory[	1045	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1046	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1047	] =	{1'b0, 6'd38, 6'd3, 3'd3};	// Note: 4A#Bb
	assign memory[	1048	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1049	] =	{1'b0, 6'd38, 6'd6, 3'd5};	// Note: 4A#Bb
	assign memory[	1050	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1051	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1052	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1053	] =	{1'b0, 6'd22, 6'd24, 3'd4};	// Note: 2F#Gb
	assign memory[	1054	] =	{1'b0, 6'd34, 6'd3, 3'd5};	// Note: 3F#Gb
	assign memory[	1055	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1056	] =	{1'b0, 6'd29, 6'd9, 3'd5};	// Note: 3C#Db
	assign memory[	1057	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1058	] =	{1'b0, 6'd29, 6'd12, 3'd3};	// Note: 3C#Db
	assign memory[	1059	] =	{1'b1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	1060	] =	{1'b0, 6'd20, 6'd18, 3'd4};	// Note: 2E
	assign memory[	1061	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1062	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1063	] =	{1'b0, 6'd39, 6'd9, 3'd3};	// Note: 4B
	assign memory[	1064	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1065	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1066	] =	{1'b0, 6'd20, 6'd6, 3'd4};	// Note: 2E
	assign memory[	1067	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1068	] =	{1'b0, 6'd20, 6'd18, 3'd4};	// Note: 2E
	assign memory[	1069	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1070	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1071	] =	{1'b0, 6'd32, 6'd9, 3'd5};	// Note: 3E
	assign memory[	1072	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1073	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1074	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1075	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1076	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1077	] =	{1'b0, 6'd17, 6'd18, 3'd4};	// Note: 2C#Db
	assign memory[	1078	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1079	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1080	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1081	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1082	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1083	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1084	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1085	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1086	] =	{1'b0, 6'd17, 6'd18, 3'd4};	// Note: 2C#Db
	assign memory[	1087	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1088	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1089	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1090	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1091	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1092	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1093	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1094	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1095	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1096	] =	{1'b0, 6'd22, 6'd6, 3'd7};	// Note: 2F#Gb
	assign memory[	1097	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1098	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1099	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1100	] =	{1'b0, 6'd24, 6'd18, 3'd7};	// Note: 2G#Ab
	assign memory[	1101	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1102	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1103	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1104	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1105	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1106	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1107	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1108	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1109	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1110	] =	{1'b0, 6'd36, 6'd24, 3'd7};	// Note: 3G#Ab
	assign memory[	1111	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1112	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1113	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1114	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1115	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1116	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1117	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1118	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1119	] =	{1'b0, 6'd30, 6'd9, 3'd5};	// Note: 3D
	assign memory[	1120	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1121	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1122	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1123	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1124	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1125	] =	{1'b0, 6'd34, 6'd24, 3'd7};	// Note: 3F#Gb
	assign memory[	1126	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1127	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1128	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1129	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1130	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1131	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1132	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1133	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1134	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1135	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1136	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1137	] =	{1'b0, 6'd38, 6'd6, 3'd5};	// Note: 4A#Bb
	assign memory[	1138	] =	{1'b0, 6'd38, 6'd12, 3'd7};	// Note: 4A#Bb
	assign memory[	1139	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1140	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1141	] =	{1'b0, 6'd34, 6'd3, 3'd5};	// Note: 3F#Gb
	assign memory[	1142	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1143	] =	{1'b0, 6'd29, 6'd6, 3'd5};	// Note: 3C#Db
	assign memory[	1144	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1145	] =	{1'b0, 6'd39, 6'd6, 3'd7};	// Note: 4B
	assign memory[	1146	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1147	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1148	] =	{1'b0, 6'd34, 6'd9, 3'd5};	// Note: 3F#Gb
	assign memory[	1149	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1150	] =	{1'b0, 6'd38, 6'd6, 3'd7};	// Note: 4A#Bb
	assign memory[	1151	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1152	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1153	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1154	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1155	] =	{1'b0, 6'd39, 6'd6, 3'd7};	// Note: 4B
	assign memory[	1156	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1157	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1158	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1159	] =	{1'b0, 6'd34, 6'd3, 3'd7};	// Note: 3F#Gb
	assign memory[	1160	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1161	] =	{1'b0, 6'd31, 6'd6, 3'd7};	// Note: 3D#Eb
	assign memory[	1162	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1163	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1164	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1165	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1166	] =	{1'b0, 6'd31, 6'd9, 3'd7};	// Note: 3D#Eb
	assign memory[	1167	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1168	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1169	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1170	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1171	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1172	] =	{1'b0, 6'd34, 6'd6, 3'd7};	// Note: 3F#Gb
	assign memory[	1173	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1174	] =	{1'b0, 6'd34, 6'd24, 3'd7};	// Note: 3F#Gb
	assign memory[	1175	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1176	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1177	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1178	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1179	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1180	] =	{1'b0, 6'd32, 6'd9, 3'd5};	// Note: 3E
	assign memory[	1181	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1182	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1183	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1184	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1185	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1186	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1187	] =	{1'b0, 6'd34, 6'd12, 3'd7};	// Note: 3F#Gb
	assign memory[	1188	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1189	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1190	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1191	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1192	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1193	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1194	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1195	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1196	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1197	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1198	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1199	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1200	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1201	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1202	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1203	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1204	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1205	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1206	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1207	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1208	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1209	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1210	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1211	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1212	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1213	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1214	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1215	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1216	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1217	] =	{1'b0, 6'd22, 6'd6, 3'd7};	// Note: 2F#Gb
	assign memory[	1218	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1219	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1220	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1221	] =	{1'b0, 6'd24, 6'd18, 3'd7};	// Note: 2G#Ab
	assign memory[	1222	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1223	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1224	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1225	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1226	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1227	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1228	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1229	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1230	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1231	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1232	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1233	] =	{1'b0, 6'd36, 6'd12, 3'd7};	// Note: 3G#Ab
	assign memory[	1234	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1235	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1236	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1237	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1238	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1239	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1240	] =	{1'b0, 6'd34, 6'd18, 3'd7};	// Note: 3F#Gb
	assign memory[	1241	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1242	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1243	] =	{1'b0, 6'd31, 6'd9, 3'd5};	// Note: 3D#Eb
	assign memory[	1244	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1245	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1246	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1247	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1248	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1249	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1250	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1251	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1252	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1253	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1254	] =	{1'b0, 6'd27, 6'd6, 3'd7};	// Note: 3B
	assign memory[	1255	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1256	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1257	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1258	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1259	] =	{1'b0, 6'd38, 6'd6, 3'd7};	// Note: 4A#Bb
	assign memory[	1260	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1261	] =	{1'b0, 6'd38, 6'd12, 3'd7};	// Note: 4A#Bb
	assign memory[	1262	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1263	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1264	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1265	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1266	] =	{1'b0, 6'd34, 6'd3, 3'd5};	// Note: 3F#Gb
	assign memory[	1267	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1268	] =	{1'b0, 6'd29, 6'd6, 3'd5};	// Note: 3C#Db
	assign memory[	1269	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1270	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1271	] =	{1'b0, 6'd34, 6'd6, 3'd7};	// Note: 3F#Gb
	assign memory[	1272	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1273	] =	{1'b0, 6'd34, 6'd9, 3'd5};	// Note: 3F#Gb
	assign memory[	1274	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1275	] =	{1'b0, 6'd34, 6'd12, 3'd7};	// Note: 3F#Gb
	assign memory[	1276	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1277	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1278	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1279	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1280	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1281	] =	{1'b0, 6'd31, 6'd6, 3'd7};	// Note: 3D#Eb
	assign memory[	1282	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1283	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1284	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1285	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1286	] =	{1'b0, 6'd29, 6'd6, 3'd7};	// Note: 3C#Db
	assign memory[	1287	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1288	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1289	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1290	] =	{1'b0, 6'd27, 6'd6, 3'd7};	// Note: 3B
	assign memory[	1291	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1292	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1293	] =	{1'b0, 6'd29, 6'd24, 3'd7};	// Note: 3C#Db
	assign memory[	1294	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1295	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1296	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1297	] =	{1'b0, 6'd29, 6'd9, 3'd5};	// Note: 3C#Db
	assign memory[	1298	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1299	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1300	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1301	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1302	] =	{1'b0, 6'd32, 6'd9, 3'd5};	// Note: 3E
	assign memory[	1303	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1304	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1305	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1306	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1307	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1308	] =	{1'b0, 6'd31, 6'd6, 3'd7};	// Note: 3D#Eb
	assign memory[	1309	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1310	] =	{1'b0, 6'd31, 6'd24, 3'd7};	// Note: 3D#Eb
	assign memory[	1311	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1312	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1313	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1314	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1315	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1316	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1317	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1318	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1319	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1320	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1321	] =	{1'b0, 6'd31, 6'd6, 3'd5};	// Note: 3D#Eb
	assign memory[	1322	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1323	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1324	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1325	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1326	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1327	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1328	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1329	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1330	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1331	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1332	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1333	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1334	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1335	] =	{1'b0, 6'd31, 6'd6, 3'd7};	// Note: 3D#Eb
	assign memory[	1336	] =	{1'b0, 6'd31, 6'd6, 3'd5};	// Note: 3D#Eb
	assign memory[	1337	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1338	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1339	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1340	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1341	] =	{1'b0, 6'd36, 6'd6, 3'd7};	// Note: 3G#Ab
	assign memory[	1342	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1343	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1344	] =	{1'b0, 6'd24, 6'd18, 3'd4};	// Note: 2G#Ab
	assign memory[	1345	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1346	] =	{1'b0, 6'd39, 6'd3, 3'd3};	// Note: 4B
	assign memory[	1347	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1348	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1349	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1350	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1351	] =	{1'b0, 6'd24, 6'd6, 3'd4};	// Note: 2G#Ab
	assign memory[	1352	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1353	] =	{1'b0, 6'd24, 6'd18, 3'd4};	// Note: 2G#Ab
	assign memory[	1354	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1355	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1356	] =	{1'b0, 6'd31, 6'd3, 3'd3};	// Note: 3D#Eb
	assign memory[	1357	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1358	] =	{1'b0, 6'd31, 6'd6, 3'd5};	// Note: 3D#Eb
	assign memory[	1359	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1360	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1361	] =	{1'b0, 6'd24, 6'd6, 3'd4};	// Note: 2G#Ab
	assign memory[	1362	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1363	] =	{1'b0, 6'd22, 6'd24, 3'd4};	// Note: 2F#Gb
	assign memory[	1364	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1365	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1366	] =	{1'b0, 6'd38, 6'd3, 3'd3};	// Note: 4A#Bb
	assign memory[	1367	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1368	] =	{1'b0, 6'd38, 6'd6, 3'd5};	// Note: 4A#Bb
	assign memory[	1369	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1370	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1371	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1372	] =	{1'b0, 6'd22, 6'd24, 3'd4};	// Note: 2F#Gb
	assign memory[	1373	] =	{1'b0, 6'd34, 6'd3, 3'd5};	// Note: 3F#Gb
	assign memory[	1374	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1375	] =	{1'b0, 6'd29, 6'd9, 3'd5};	// Note: 3C#Db
	assign memory[	1376	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1377	] =	{1'b0, 6'd29, 6'd12, 3'd3};	// Note: 3C#Db
	assign memory[	1378	] =	{1'b1, 6'd0, 6'd12, 3'd0};	// Note: rest
	assign memory[	1379	] =	{1'b0, 6'd20, 6'd18, 3'd4};	// Note: 2E
	assign memory[	1380	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1381	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1382	] =	{1'b0, 6'd39, 6'd9, 3'd3};	// Note: 4B
	assign memory[	1383	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1384	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1385	] =	{1'b0, 6'd20, 6'd6, 3'd4};	// Note: 2E
	assign memory[	1386	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1387	] =	{1'b0, 6'd20, 6'd18, 3'd4};	// Note: 2E
	assign memory[	1388	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1389	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1390	] =	{1'b0, 6'd32, 6'd9, 3'd5};	// Note: 3E
	assign memory[	1391	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1392	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1393	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1394	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1395	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1396	] =	{1'b0, 6'd17, 6'd18, 3'd4};	// Note: 2C#Db
	assign memory[	1397	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1398	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1399	] =	{1'b1, 6'd0, 6'd9, 3'd0};	// Note: rest
	assign memory[	1400	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1401	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1402	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1403	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1404	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1405	] =	{1'b0, 6'd17, 6'd18, 3'd4};	// Note: 2C#Db
	assign memory[	1406	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1407	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1408	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1409	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1410	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1411	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1412	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1413	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1414	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1415	] =	{1'b0, 6'd22, 6'd6, 3'd7};	// Note: 2F#Gb
	assign memory[	1416	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1417	] =	{1'b0, 6'd17, 6'd6, 3'd4};	// Note: 2C#Db
	assign memory[	1418	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1419	] =	{1'b0, 6'd24, 6'd18, 3'd7};	// Note: 2G#Ab
	assign memory[	1420	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1421	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1422	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1423	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1424	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1425	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1426	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1427	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1428	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1429	] =	{1'b0, 6'd36, 6'd24, 3'd7};	// Note: 3G#Ab
	assign memory[	1430	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1431	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1432	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1433	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1434	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1435	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1436	] =	{1'b0, 6'd12, 6'd6, 3'd3};	// Note: 1G#Ab
	assign memory[	1437	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1438	] =	{1'b0, 6'd30, 6'd9, 3'd5};	// Note: 3D
	assign memory[	1439	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1440	] =	{1'b0, 6'd12, 6'd6, 3'd4};	// Note: 1G#Ab
	assign memory[	1441	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1442	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1443	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1444	] =	{1'b0, 6'd34, 6'd24, 3'd7};	// Note: 3F#Gb
	assign memory[	1445	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1446	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1447	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1448	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1449	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1450	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1451	] =	{1'b0, 6'd38, 6'd9, 3'd5};	// Note: 4A#Bb
	assign memory[	1452	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1453	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1454	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1455	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1456	] =	{1'b0, 6'd38, 6'd6, 3'd5};	// Note: 4A#Bb
	assign memory[	1457	] =	{1'b0, 6'd38, 6'd12, 3'd7};	// Note: 4A#Bb
	assign memory[	1458	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1459	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1460	] =	{1'b0, 6'd34, 6'd3, 3'd5};	// Note: 3F#Gb
	assign memory[	1461	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1462	] =	{1'b0, 6'd29, 6'd6, 3'd5};	// Note: 3C#Db
	assign memory[	1463	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1464	] =	{1'b0, 6'd39, 6'd6, 3'd7};	// Note: 4B
	assign memory[	1465	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1466	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1467	] =	{1'b0, 6'd34, 6'd9, 3'd5};	// Note: 3F#Gb
	assign memory[	1468	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1469	] =	{1'b0, 6'd38, 6'd6, 3'd7};	// Note: 4A#Bb
	assign memory[	1470	] =	{1'b0, 6'd10, 6'd6, 3'd4};	// Note: 1F#Gb
	assign memory[	1471	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1472	] =	{1'b0, 6'd10, 6'd6, 3'd3};	// Note: 1F#Gb
	assign memory[	1473	] =	{1'b0, 6'd34, 6'd6, 3'd5};	// Note: 3F#Gb
	assign memory[	1474	] =	{1'b0, 6'd39, 6'd6, 3'd7};	// Note: 4B
	assign memory[	1475	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1476	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1477	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1478	] =	{1'b0, 6'd34, 6'd3, 3'd7};	// Note: 3F#Gb
	assign memory[	1479	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1480	] =	{1'b0, 6'd31, 6'd6, 3'd7};	// Note: 3D#Eb
	assign memory[	1481	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1482	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1483	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1484	] =	{1'b0, 6'd39, 6'd9, 3'd5};	// Note: 4B
	assign memory[	1485	] =	{1'b0, 6'd31, 6'd9, 3'd7};	// Note: 3D#Eb
	assign memory[	1486	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1487	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1488	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1489	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1490	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1491	] =	{1'b0, 6'd34, 6'd6, 3'd7};	// Note: 3F#Gb
	assign memory[	1492	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1493	] =	{1'b0, 6'd34, 6'd24, 3'd7};	// Note: 3F#Gb
	assign memory[	1494	] =	{1'b0, 6'd36, 6'd9, 3'd5};	// Note: 3G#Ab
	assign memory[	1495	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1496	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1497	] =	{1'b0, 6'd8, 6'd6, 3'd3};	// Note: 1E
	assign memory[	1498	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1499	] =	{1'b0, 6'd32, 6'd9, 3'd5};	// Note: 3E
	assign memory[	1500	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1501	] =	{1'b0, 6'd8, 6'd6, 3'd4};	// Note: 1E
	assign memory[	1502	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1503	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1504	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1505	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1506	] =	{1'b0, 6'd34, 6'd12, 3'd7};	// Note: 3F#Gb
	assign memory[	1507	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1508	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1509	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1510	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1511	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1512	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1513	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1514	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1515	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1516	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1517	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1518	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1519	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1520	] =	{1'b0, 6'd39, 6'd6, 3'd5};	// Note: 4B
	assign memory[	1521	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest
	assign memory[	1522	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1523	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1524	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1525	] =	{1'b0, 6'd36, 6'd6, 3'd5};	// Note: 3G#Ab
	assign memory[	1526	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1527	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1528	] =	{1'b0, 6'd5, 6'd6, 3'd3};	// Note: 1C#Db
	assign memory[	1529	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1530	] =	{1'b0, 6'd39, 6'd3, 3'd5};	// Note: 4B
	assign memory[	1531	] =	{1'b1, 6'd0, 6'd3, 3'd0};	// Note: rest
	assign memory[	1532	] =	{1'b0, 6'd24, 6'd6, 3'd7};	// Note: 2G#Ab
	assign memory[	1533	] =	{1'b0, 6'd32, 6'd6, 3'd5};	// Note: 3E
	assign memory[	1534	] =	{1'b0, 6'd5, 6'd6, 3'd4};	// Note: 1C#Db
	assign memory[	1535	] =	{1'b1, 6'd0, 6'd6, 3'd0};	// Note: rest

// Song 4

	assign memory[	1536	] =	{1'b0, 6'd26, 6'd48, 3'd3};	// Note: 3A#Bb
	assign memory[	1537	] =	{1'b0, 6'd33, 6'd48, 3'd3};	// Note: 3F
	assign memory[	1538	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1539	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1540	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1541	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1542	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1543	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1544	] =	{1'b0, 6'd49, 6'd8, 3'd4};	// Note: 5A
	assign memory[	1545	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1546	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1547	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1548	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1549	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1550	] =	{1'b0, 6'd26, 6'd48, 3'd3};	// Note: 3A#Bb
	assign memory[	1551	] =	{1'b0, 6'd33, 6'd48, 3'd3};	// Note: 3F
	assign memory[	1552	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1553	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1554	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1555	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1556	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1557	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1558	] =	{1'b0, 6'd49, 6'd8, 3'd4};	// Note: 5A
	assign memory[	1559	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1560	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1561	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1562	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1563	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1564	] =	{1'b0, 6'd23, 6'd48, 3'd4};	// Note: 2G
	assign memory[	1565	] =	{1'b0, 6'd30, 6'd48, 3'd4};	// Note: 3D
	assign memory[	1566	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1567	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1568	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1569	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1570	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1571	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1572	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1573	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1574	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1575	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1576	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1577	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1578	] =	{1'b0, 6'd23, 6'd48, 3'd4};	// Note: 2G
	assign memory[	1579	] =	{1'b0, 6'd30, 6'd48, 3'd4};	// Note: 3D
	assign memory[	1580	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1581	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1582	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1583	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1584	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1585	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1586	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1587	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1588	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1589	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1590	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1591	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1592	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1593	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1594	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1595	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1596	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1597	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1598	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1599	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1600	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1601	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1602	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1603	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1604	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1605	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1606	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1607	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1608	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1609	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1610	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1611	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1612	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1613	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1614	] =	{1'b0, 6'd44, 6'd8, 3'd4};	// Note: 4E
	assign memory[	1615	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1616	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1617	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1618	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1619	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1620	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1621	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1622	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1623	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1624	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1625	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1626	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1627	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1628	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1629	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1630	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1631	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1632	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1633	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1634	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1635	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1636	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1637	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1638	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1639	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1640	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1641	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1642	] =	{1'b0, 6'd44, 6'd8, 3'd4};	// Note: 4E
	assign memory[	1643	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1644	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1645	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1646	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1647	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1648	] =	{1'b0, 6'd26, 6'd48, 3'd3};	// Note: 3A#Bb
	assign memory[	1649	] =	{1'b0, 6'd33, 6'd48, 3'd3};	// Note: 3F
	assign memory[	1650	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1651	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1652	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1653	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1654	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1655	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1656	] =	{1'b0, 6'd49, 6'd8, 3'd4};	// Note: 5A
	assign memory[	1657	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1658	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1659	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1660	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1661	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1662	] =	{1'b0, 6'd26, 6'd48, 3'd3};	// Note: 3A#Bb
	assign memory[	1663	] =	{1'b0, 6'd33, 6'd48, 3'd3};	// Note: 3F
	assign memory[	1664	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1665	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1666	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1667	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1668	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1669	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1670	] =	{1'b0, 6'd49, 6'd8, 3'd4};	// Note: 5A
	assign memory[	1671	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1672	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1673	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1674	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1675	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1676	] =	{1'b0, 6'd23, 6'd48, 3'd4};	// Note: 2G
	assign memory[	1677	] =	{1'b0, 6'd30, 6'd48, 3'd4};	// Note: 3D
	assign memory[	1678	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1679	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1680	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1681	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1682	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1683	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1684	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1685	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1686	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1687	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1688	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1689	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1690	] =	{1'b0, 6'd23, 6'd48, 3'd4};	// Note: 2G
	assign memory[	1691	] =	{1'b0, 6'd30, 6'd48, 3'd4};	// Note: 3D
	assign memory[	1692	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1693	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1694	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1695	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1696	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1697	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1698	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1699	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1700	] =	{1'b0, 6'd38, 6'd8, 3'd4};	// Note: 4A#Bb
	assign memory[	1701	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1702	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1703	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1704	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1705	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1706	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1707	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1708	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1709	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1710	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1711	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1712	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1713	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1714	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1715	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1716	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1717	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1718	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1719	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1720	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1721	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1722	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1723	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1724	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1725	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1726	] =	{1'b0, 6'd44, 6'd8, 3'd4};	// Note: 4E
	assign memory[	1727	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1728	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1729	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1730	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1731	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1732	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1733	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1734	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1735	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1736	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1737	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1738	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1739	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1740	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1741	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1742	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1743	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1744	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1745	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1746	] =	{1'b0, 6'd18, 6'd48, 3'd3};	// Note: 2D
	assign memory[	1747	] =	{1'b0, 6'd30, 6'd48, 3'd3};	// Note: 3D
	assign memory[	1748	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1749	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1750	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1751	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1752	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1753	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1754	] =	{1'b0, 6'd44, 6'd8, 3'd4};	// Note: 4E
	assign memory[	1755	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1756	] =	{1'b0, 6'd37, 6'd8, 3'd4};	// Note: 4A
	assign memory[	1757	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1758	] =	{1'b0, 6'd45, 6'd8, 3'd4};	// Note: 4F
	assign memory[	1759	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1760	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1761	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1762	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1763	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1764	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1765	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1766	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1767	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1768	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1769	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1770	] =	{1'b0, 6'd49, 6'd8, 3'd7};	// Note: 5
	assign memory[	1771	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1772	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1773	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1774	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1775	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1776	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1777	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1778	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1779	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1780	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1781	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1782	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1783	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1784	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1785	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1786	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1787	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1788	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1789	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1790	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1791	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1792	] =	{1'b0, 6'd49, 6'd8, 3'd7};	// Note: 5A
	assign memory[	1793	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1794	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1795	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1796	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1797	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1798	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1799	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1800	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1801	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1802	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1803	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1804	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1805	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1806	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1807	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1808	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1809	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1810	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1811	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1812	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1813	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1814	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1815	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1816	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1817	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1818	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1819	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1820	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1821	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1822	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1823	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1824	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1825	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1826	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1827	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1828	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1829	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1830	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1831	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1832	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1833	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1834	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1835	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1836	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1837	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1838	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1839	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1840	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1841	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1842	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1843	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1844	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1845	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1846	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1847	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1848	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1849	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1850	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1851	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1852	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1853	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1854	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1855	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1856	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1857	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1858	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1859	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1860	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1861	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1862	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1863	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1864	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1865	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1866	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1867	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1868	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1869	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1870	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1871	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1872	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1873	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1874	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1875	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1876	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1877	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1878	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1879	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1880	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1881	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1882	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1883	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1884	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1885	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1886	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1887	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1888	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1889	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1890	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1891	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1892	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1893	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1894	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1895	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1896	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1897	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1898	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1899	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1900	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1901	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1902	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1903	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1904	] =	{1'b0, 6'd46, 6'd8, 3'd6};	// Note: 4F#Gb
	assign memory[	1905	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1906	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1907	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1908	] =	{1'b0, 6'd46, 6'd8, 3'd3};	// Note: 4F#Gb
	assign memory[	1909	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1910	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1911	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1912	] =	{1'b0, 6'd46, 6'd8, 3'd3};	// Note: 4F#Gb
	assign memory[	1913	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1914	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1915	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1916	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1917	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	1918	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1919	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1920	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1921	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1922	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	1923	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1924	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1925	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	1926	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1927	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1928	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1929	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1930	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1931	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1932	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1933	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1934	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1935	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1936	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1937	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1938	] =	{1'b0, 6'd49, 6'd8, 3'd7};	// Note: 5A
	assign memory[	1939	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1940	] =	{1'b0, 6'd26, 6'd8, 3'd6};	// Note: 3A#Bb
	assign memory[	1941	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1942	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1943	] =	{1'b0, 6'd26, 6'd8, 3'd3};	// Note: 3A#Bb
	assign memory[	1944	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1945	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1946	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1947	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1948	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1949	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1950	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1951	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1952	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1953	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1954	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1955	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1956	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1957	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1958	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1959	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1960	] =	{1'b0, 6'd49, 6'd8, 3'd7};	// Note: 5A
	assign memory[	1961	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1962	] =	{1'b0, 6'd33, 6'd8, 3'd6};	// Note: 3F
	assign memory[	1963	] =	{1'b0, 6'd37, 6'd8, 3'd6};	// Note: 4A
	assign memory[	1964	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1965	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1966	] =	{1'b0, 6'd33, 6'd8, 3'd3};	// Note: 3F
	assign memory[	1967	] =	{1'b0, 6'd37, 6'd8, 3'd3};	// Note: 4A
	assign memory[	1968	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1969	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1970	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1971	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1972	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1973	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1974	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1975	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1976	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1977	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1978	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1979	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1980	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	1981	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1982	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1983	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1984	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1985	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1986	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	1987	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1988	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1989	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1990	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1991	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1992	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	1993	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	1994	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	1995	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	1996	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	1997	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	1998	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	1999	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2000	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	2001	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	2002	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	2003	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2004	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	2005	] =	{1'b0, 6'd23, 6'd8, 3'd6};	// Note: 2G
	assign memory[	2006	] =	{1'b0, 6'd38, 6'd8, 3'd7};	// Note: 4A#Bb
	assign memory[	2007	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2008	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	2009	] =	{1'b0, 6'd23, 6'd8, 3'd3};	// Note: 2G
	assign memory[	2010	] =	{1'b0, 6'd40, 6'd8, 3'd4};	// Note: 4C
	assign memory[	2011	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2012	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	2013	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	2014	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2015	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	2016	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	2017	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2018	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	2019	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	2020	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2021	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	2022	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	2023	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2024	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	2025	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	2026	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2027	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	2028	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	2029	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2030	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	2031	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	2032	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	2033	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2034	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	2035	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	2036	] =	{1'b0, 6'd40, 6'd8, 3'd7};	// Note: 4C
	assign memory[	2037	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2038	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	2039	] =	{1'b0, 6'd18, 6'd8, 3'd6};	// Note: 2D
	assign memory[	2040	] =	{1'b0, 6'd37, 6'd8, 3'd7};	// Note: 4A
	assign memory[	2041	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2042	] =	{1'b0, 6'd47, 6'd8, 3'd3};	// Note: 4G
	assign memory[	2043	] =	{1'b0, 6'd18, 6'd8, 3'd3};	// Note: 2D
	assign memory[	2044	] =	{1'b0, 6'd45, 6'd8, 3'd7};	// Note: 4F
	assign memory[	2045	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
	assign memory[	2046	] =	{1'b0, 6'd47, 6'd8, 3'd6};	// Note: 4G
	assign memory[	2047	] =	{1'b1, 6'd0, 6'd8, 3'd0};	// Note: rest
					
endmodule