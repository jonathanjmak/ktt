
    );


endmodule
